library ieee;

use ieee.std_logic_1164.all;

entity pixelGenerator_tb is

end pixelGenerator_tb;

architecture structural of pixelGenerator_tb is
	component
begin

end structrual;
