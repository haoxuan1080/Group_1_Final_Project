library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pixelGenerator is
	port(
			clk, ROM_clk, rst_n, video_on, eof 				: in std_logic;
			xx , yy, x_b, y_b													: in natural;
			pixel_row, pixel_column						    : in std_logic_vector(9 downto 0);
		
			red_out, green_out, blue_out					: out std_logic_vector(7 downto 0)
		);
end entity pixelGenerator;

architecture behavioral of pixelGenerator is

constant color_red 	 	 : std_logic_vector(2 downto 0) := "000";
constant color_green	 : std_logic_vector(2 downto 0) := "001";
constant color_blue 	 : std_logic_vector(2 downto 0) := "010";
constant color_yellow 	 : std_logic_vector(2 downto 0) := "011";
constant color_magenta 	 : std_logic_vector(2 downto 0) := "100";
constant color_cyan 	 : std_logic_vector(2 downto 0) := "101";
constant color_black 	 : std_logic_vector(2 downto 0) := "110";
constant color_white	 : std_logic_vector(2 downto 0) := "111";
	
component colorDecoder is
	port
	(
		address		: in std_logic_vector (2 downto 0);
		q			: out std_logic_vector (23 downto 0)
	);
end component colorDecoder;

signal pixel_row_int, pixel_column_int 				: natural;
signal colorAddress : std_logic_vector (2 downto 0);
signal color        : std_logic_vector (23 downto 0);

begin
--------------------------------------------------------------------------------------------
	
	red_out <= color(23 downto 16);
	green_out <= color(15 downto 8);
	blue_out <= color(7 downto 0);

	pixel_row_int <= to_integer(unsigned(pixel_row));
	pixel_column_int <= to_integer(unsigned(pixel_column));
	
--------------------------------------------------------------------------------------------	
	colors : colorDecoder
		port map(colorAddress,color);
--------------------------------------------------------------------------------------------	

	pixelDraw : process(clk, rst_n) is
	
	begin
	
		if (rst_n = '0')then
			colorAddress <= color_white; 			
		elsif (rising_edge(clk)) then
			if ((abs(pixel_row_int - xx) < 10) and (abs(pixel_column_int -yy) < 5)) then
				colorAddress <= color_yellow;
			elsif((abs(pixel_row_int - x_b) < 5) and (abs(pixel_column_int -y_b) < 2))then
				colorAddress <= color_blue;
			else
				colorAddress <= color_cyan;
			end if;
			
		end if;
		
	end process pixelDraw;	

--------------------------------------------------------------------------------------------
	
end architecture behavioral;		