library ieee;

use ieee.std_logic_1164.all;
	
package Game_constant is
	constant Screen_Width: natural :=640;
	constant Screen_Height: natural :=480;
	constant Tank_Width: natural:=30;
	constant Tank_Hight: natural:=20;

	constant Bullet_Radius: natural:=5;

end package Game_constant;

package body Game_constant is

end package body Game_constant;
